module sing(
    input [9:0] P1X;
    input [9:0] P1Y;

    input [9:0] P2X;
    input [9:0] P2Y;

    input [9:0] PTX;
    input [9:0] PTY;
);

    wire 
